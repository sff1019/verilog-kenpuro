module target_square();
  wire [11:0] w_sq_pos_x, w_sq_pos_y;

  
